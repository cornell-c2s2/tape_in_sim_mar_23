
`ifndef FFT_VRTL
`define FFT_VRTL

`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/TwiddleGeneratorVRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_512VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_256VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_128VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_64VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_32VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_16VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_8VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_2VRTL.v"
`include "../FFT/FFT-Twiddle_Generator/sim/FFTTwiddleGenerator/SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_4VRTL.v"
`include "../FFT/FFT-Crossbar/sim/CombinationalFFTCrossbar/CombinationalFFTCrossbarVRTL.v"
`include "../FFT/FFT_StageVRTL.v"
module FFTVRTL 
   #(
        BIT_WIDTH  = 32,
        DECIMAL_PT = 16,
        N_SAMPLES  = 8
    )
    (
        input  logic [BIT_WIDTH - 1:0] recv_msg [N_SAMPLES - 1:0],
        input  logic                   recv_val                  ,
        output logic                   recv_rdy                  ,

        output logic [BIT_WIDTH - 1:0] send_msg [N_SAMPLES - 1:0],
        output logic                   send_val                  ,
        input  logic                   send_rdy                  ,

        input  logic                   reset                     ,
        input  logic                   clk
    );

    logic [BIT_WIDTH - 1:0] real_msg       [$clog2(N_SAMPLES):0][N_SAMPLES - 1:0];
    logic [BIT_WIDTH - 1:0] complex_msg    [$clog2(N_SAMPLES):0][N_SAMPLES - 1:0];

    logic                   val_in         [$clog2(N_SAMPLES):0];
    logic                   rdy_in         [$clog2(N_SAMPLES):0];

    logic [BIT_WIDTH - 1:0] sine_wave_out [0:N_SAMPLES - 1];


    assign val_in  [0] = recv_val;
    assign recv_rdy    = rdy_in[0];

    assign send_val                  = val_in     [$clog2(N_SAMPLES)];
    assign rdy_in[$clog2(N_SAMPLES)] = send_rdy;

    


    always @(*) begin
        int i;
        for(i = 0; i < N_SAMPLES; i++) begin
            complex_msg[0][i] = 0;
        end
    end

    //Manual 8-bit bit reversal TODO make parametrized
    generate
        if(N_SAMPLES == 512) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][256] = recv_msg[1];
            assign real_msg[0][128] = recv_msg[2];
            assign real_msg[0][384] = recv_msg[3];
            assign real_msg[0][64] = recv_msg[4];
            assign real_msg[0][320] = recv_msg[5];
            assign real_msg[0][192] = recv_msg[6];
            assign real_msg[0][448] = recv_msg[7];
            assign real_msg[0][32] = recv_msg[8];
            assign real_msg[0][288] = recv_msg[9];
            assign real_msg[0][160] = recv_msg[10];
            assign real_msg[0][416] = recv_msg[11];
            assign real_msg[0][96] = recv_msg[12];
            assign real_msg[0][352] = recv_msg[13];
            assign real_msg[0][224] = recv_msg[14];
            assign real_msg[0][480] = recv_msg[15];
            assign real_msg[0][16] = recv_msg[16];
            assign real_msg[0][272] = recv_msg[17];
            assign real_msg[0][144] = recv_msg[18];
            assign real_msg[0][400] = recv_msg[19];
            assign real_msg[0][80] = recv_msg[20];
            assign real_msg[0][336] = recv_msg[21];
            assign real_msg[0][208] = recv_msg[22];
            assign real_msg[0][464] = recv_msg[23];
            assign real_msg[0][48] = recv_msg[24];
            assign real_msg[0][304] = recv_msg[25];
            assign real_msg[0][176] = recv_msg[26];
            assign real_msg[0][432] = recv_msg[27];
            assign real_msg[0][112] = recv_msg[28];
            assign real_msg[0][368] = recv_msg[29];
            assign real_msg[0][240] = recv_msg[30];
            assign real_msg[0][496] = recv_msg[31];
            assign real_msg[0][8] = recv_msg[32];
            assign real_msg[0][264] = recv_msg[33];
            assign real_msg[0][136] = recv_msg[34];
            assign real_msg[0][392] = recv_msg[35];
            assign real_msg[0][72] = recv_msg[36];
            assign real_msg[0][328] = recv_msg[37];
            assign real_msg[0][200] = recv_msg[38];
            assign real_msg[0][456] = recv_msg[39];
            assign real_msg[0][40] = recv_msg[40];
            assign real_msg[0][296] = recv_msg[41];
            assign real_msg[0][168] = recv_msg[42];
            assign real_msg[0][424] = recv_msg[43];
            assign real_msg[0][104] = recv_msg[44];
            assign real_msg[0][360] = recv_msg[45];
            assign real_msg[0][232] = recv_msg[46];
            assign real_msg[0][488] = recv_msg[47];
            assign real_msg[0][24] = recv_msg[48];
            assign real_msg[0][280] = recv_msg[49];
            assign real_msg[0][152] = recv_msg[50];
            assign real_msg[0][408] = recv_msg[51];
            assign real_msg[0][88] = recv_msg[52];
            assign real_msg[0][344] = recv_msg[53];
            assign real_msg[0][216] = recv_msg[54];
            assign real_msg[0][472] = recv_msg[55];
            assign real_msg[0][56] = recv_msg[56];
            assign real_msg[0][312] = recv_msg[57];
            assign real_msg[0][184] = recv_msg[58];
            assign real_msg[0][440] = recv_msg[59];
            assign real_msg[0][120] = recv_msg[60];
            assign real_msg[0][376] = recv_msg[61];
            assign real_msg[0][248] = recv_msg[62];
            assign real_msg[0][504] = recv_msg[63];
            assign real_msg[0][4] = recv_msg[64];
            assign real_msg[0][260] = recv_msg[65];
            assign real_msg[0][132] = recv_msg[66];
            assign real_msg[0][388] = recv_msg[67];
            assign real_msg[0][68] = recv_msg[68];
            assign real_msg[0][324] = recv_msg[69];
            assign real_msg[0][196] = recv_msg[70];
            assign real_msg[0][452] = recv_msg[71];
            assign real_msg[0][36] = recv_msg[72];
            assign real_msg[0][292] = recv_msg[73];
            assign real_msg[0][164] = recv_msg[74];
            assign real_msg[0][420] = recv_msg[75];
            assign real_msg[0][100] = recv_msg[76];
            assign real_msg[0][356] = recv_msg[77];
            assign real_msg[0][228] = recv_msg[78];
            assign real_msg[0][484] = recv_msg[79];
            assign real_msg[0][20] = recv_msg[80];
            assign real_msg[0][276] = recv_msg[81];
            assign real_msg[0][148] = recv_msg[82];
            assign real_msg[0][404] = recv_msg[83];
            assign real_msg[0][84] = recv_msg[84];
            assign real_msg[0][340] = recv_msg[85];
            assign real_msg[0][212] = recv_msg[86];
            assign real_msg[0][468] = recv_msg[87];
            assign real_msg[0][52] = recv_msg[88];
            assign real_msg[0][308] = recv_msg[89];
            assign real_msg[0][180] = recv_msg[90];
            assign real_msg[0][436] = recv_msg[91];
            assign real_msg[0][116] = recv_msg[92];
            assign real_msg[0][372] = recv_msg[93];
            assign real_msg[0][244] = recv_msg[94];
            assign real_msg[0][500] = recv_msg[95];
            assign real_msg[0][12] = recv_msg[96];
            assign real_msg[0][268] = recv_msg[97];
            assign real_msg[0][140] = recv_msg[98];
            assign real_msg[0][396] = recv_msg[99];
            assign real_msg[0][76] = recv_msg[100];
            assign real_msg[0][332] = recv_msg[101];
            assign real_msg[0][204] = recv_msg[102];
            assign real_msg[0][460] = recv_msg[103];
            assign real_msg[0][44] = recv_msg[104];
            assign real_msg[0][300] = recv_msg[105];
            assign real_msg[0][172] = recv_msg[106];
            assign real_msg[0][428] = recv_msg[107];
            assign real_msg[0][108] = recv_msg[108];
            assign real_msg[0][364] = recv_msg[109];
            assign real_msg[0][236] = recv_msg[110];
            assign real_msg[0][492] = recv_msg[111];
            assign real_msg[0][28] = recv_msg[112];
            assign real_msg[0][284] = recv_msg[113];
            assign real_msg[0][156] = recv_msg[114];
            assign real_msg[0][412] = recv_msg[115];
            assign real_msg[0][92] = recv_msg[116];
            assign real_msg[0][348] = recv_msg[117];
            assign real_msg[0][220] = recv_msg[118];
            assign real_msg[0][476] = recv_msg[119];
            assign real_msg[0][60] = recv_msg[120];
            assign real_msg[0][316] = recv_msg[121];
            assign real_msg[0][188] = recv_msg[122];
            assign real_msg[0][444] = recv_msg[123];
            assign real_msg[0][124] = recv_msg[124];
            assign real_msg[0][380] = recv_msg[125];
            assign real_msg[0][252] = recv_msg[126];
            assign real_msg[0][508] = recv_msg[127];
            assign real_msg[0][2] = recv_msg[128];
            assign real_msg[0][258] = recv_msg[129];
            assign real_msg[0][130] = recv_msg[130];
            assign real_msg[0][386] = recv_msg[131];
            assign real_msg[0][66] = recv_msg[132];
            assign real_msg[0][322] = recv_msg[133];
            assign real_msg[0][194] = recv_msg[134];
            assign real_msg[0][450] = recv_msg[135];
            assign real_msg[0][34] = recv_msg[136];
            assign real_msg[0][290] = recv_msg[137];
            assign real_msg[0][162] = recv_msg[138];
            assign real_msg[0][418] = recv_msg[139];
            assign real_msg[0][98] = recv_msg[140];
            assign real_msg[0][354] = recv_msg[141];
            assign real_msg[0][226] = recv_msg[142];
            assign real_msg[0][482] = recv_msg[143];
            assign real_msg[0][18] = recv_msg[144];
            assign real_msg[0][274] = recv_msg[145];
            assign real_msg[0][146] = recv_msg[146];
            assign real_msg[0][402] = recv_msg[147];
            assign real_msg[0][82] = recv_msg[148];
            assign real_msg[0][338] = recv_msg[149];
            assign real_msg[0][210] = recv_msg[150];
            assign real_msg[0][466] = recv_msg[151];
            assign real_msg[0][50] = recv_msg[152];
            assign real_msg[0][306] = recv_msg[153];
            assign real_msg[0][178] = recv_msg[154];
            assign real_msg[0][434] = recv_msg[155];
            assign real_msg[0][114] = recv_msg[156];
            assign real_msg[0][370] = recv_msg[157];
            assign real_msg[0][242] = recv_msg[158];
            assign real_msg[0][498] = recv_msg[159];
            assign real_msg[0][10] = recv_msg[160];
            assign real_msg[0][266] = recv_msg[161];
            assign real_msg[0][138] = recv_msg[162];
            assign real_msg[0][394] = recv_msg[163];
            assign real_msg[0][74] = recv_msg[164];
            assign real_msg[0][330] = recv_msg[165];
            assign real_msg[0][202] = recv_msg[166];
            assign real_msg[0][458] = recv_msg[167];
            assign real_msg[0][42] = recv_msg[168];
            assign real_msg[0][298] = recv_msg[169];
            assign real_msg[0][170] = recv_msg[170];
            assign real_msg[0][426] = recv_msg[171];
            assign real_msg[0][106] = recv_msg[172];
            assign real_msg[0][362] = recv_msg[173];
            assign real_msg[0][234] = recv_msg[174];
            assign real_msg[0][490] = recv_msg[175];
            assign real_msg[0][26] = recv_msg[176];
            assign real_msg[0][282] = recv_msg[177];
            assign real_msg[0][154] = recv_msg[178];
            assign real_msg[0][410] = recv_msg[179];
            assign real_msg[0][90] = recv_msg[180];
            assign real_msg[0][346] = recv_msg[181];
            assign real_msg[0][218] = recv_msg[182];
            assign real_msg[0][474] = recv_msg[183];
            assign real_msg[0][58] = recv_msg[184];
            assign real_msg[0][314] = recv_msg[185];
            assign real_msg[0][186] = recv_msg[186];
            assign real_msg[0][442] = recv_msg[187];
            assign real_msg[0][122] = recv_msg[188];
            assign real_msg[0][378] = recv_msg[189];
            assign real_msg[0][250] = recv_msg[190];
            assign real_msg[0][506] = recv_msg[191];
            assign real_msg[0][6] = recv_msg[192];
            assign real_msg[0][262] = recv_msg[193];
            assign real_msg[0][134] = recv_msg[194];
            assign real_msg[0][390] = recv_msg[195];
            assign real_msg[0][70] = recv_msg[196];
            assign real_msg[0][326] = recv_msg[197];
            assign real_msg[0][198] = recv_msg[198];
            assign real_msg[0][454] = recv_msg[199];
            assign real_msg[0][38] = recv_msg[200];
            assign real_msg[0][294] = recv_msg[201];
            assign real_msg[0][166] = recv_msg[202];
            assign real_msg[0][422] = recv_msg[203];
            assign real_msg[0][102] = recv_msg[204];
            assign real_msg[0][358] = recv_msg[205];
            assign real_msg[0][230] = recv_msg[206];
            assign real_msg[0][486] = recv_msg[207];
            assign real_msg[0][22] = recv_msg[208];
            assign real_msg[0][278] = recv_msg[209];
            assign real_msg[0][150] = recv_msg[210];
            assign real_msg[0][406] = recv_msg[211];
            assign real_msg[0][86] = recv_msg[212];
            assign real_msg[0][342] = recv_msg[213];
            assign real_msg[0][214] = recv_msg[214];
            assign real_msg[0][470] = recv_msg[215];
            assign real_msg[0][54] = recv_msg[216];
            assign real_msg[0][310] = recv_msg[217];
            assign real_msg[0][182] = recv_msg[218];
            assign real_msg[0][438] = recv_msg[219];
            assign real_msg[0][118] = recv_msg[220];
            assign real_msg[0][374] = recv_msg[221];
            assign real_msg[0][246] = recv_msg[222];
            assign real_msg[0][502] = recv_msg[223];
            assign real_msg[0][14] = recv_msg[224];
            assign real_msg[0][270] = recv_msg[225];
            assign real_msg[0][142] = recv_msg[226];
            assign real_msg[0][398] = recv_msg[227];
            assign real_msg[0][78] = recv_msg[228];
            assign real_msg[0][334] = recv_msg[229];
            assign real_msg[0][206] = recv_msg[230];
            assign real_msg[0][462] = recv_msg[231];
            assign real_msg[0][46] = recv_msg[232];
            assign real_msg[0][302] = recv_msg[233];
            assign real_msg[0][174] = recv_msg[234];
            assign real_msg[0][430] = recv_msg[235];
            assign real_msg[0][110] = recv_msg[236];
            assign real_msg[0][366] = recv_msg[237];
            assign real_msg[0][238] = recv_msg[238];
            assign real_msg[0][494] = recv_msg[239];
            assign real_msg[0][30] = recv_msg[240];
            assign real_msg[0][286] = recv_msg[241];
            assign real_msg[0][158] = recv_msg[242];
            assign real_msg[0][414] = recv_msg[243];
            assign real_msg[0][94] = recv_msg[244];
            assign real_msg[0][350] = recv_msg[245];
            assign real_msg[0][222] = recv_msg[246];
            assign real_msg[0][478] = recv_msg[247];
            assign real_msg[0][62] = recv_msg[248];
            assign real_msg[0][318] = recv_msg[249];
            assign real_msg[0][190] = recv_msg[250];
            assign real_msg[0][446] = recv_msg[251];
            assign real_msg[0][126] = recv_msg[252];
            assign real_msg[0][382] = recv_msg[253];
            assign real_msg[0][254] = recv_msg[254];
            assign real_msg[0][510] = recv_msg[255];
            assign real_msg[0][1] = recv_msg[256];
            assign real_msg[0][257] = recv_msg[257];
            assign real_msg[0][129] = recv_msg[258];
            assign real_msg[0][385] = recv_msg[259];
            assign real_msg[0][65] = recv_msg[260];
            assign real_msg[0][321] = recv_msg[261];
            assign real_msg[0][193] = recv_msg[262];
            assign real_msg[0][449] = recv_msg[263];
            assign real_msg[0][33] = recv_msg[264];
            assign real_msg[0][289] = recv_msg[265];
            assign real_msg[0][161] = recv_msg[266];
            assign real_msg[0][417] = recv_msg[267];
            assign real_msg[0][97] = recv_msg[268];
            assign real_msg[0][353] = recv_msg[269];
            assign real_msg[0][225] = recv_msg[270];
            assign real_msg[0][481] = recv_msg[271];
            assign real_msg[0][17] = recv_msg[272];
            assign real_msg[0][273] = recv_msg[273];
            assign real_msg[0][145] = recv_msg[274];
            assign real_msg[0][401] = recv_msg[275];
            assign real_msg[0][81] = recv_msg[276];
            assign real_msg[0][337] = recv_msg[277];
            assign real_msg[0][209] = recv_msg[278];
            assign real_msg[0][465] = recv_msg[279];
            assign real_msg[0][49] = recv_msg[280];
            assign real_msg[0][305] = recv_msg[281];
            assign real_msg[0][177] = recv_msg[282];
            assign real_msg[0][433] = recv_msg[283];
            assign real_msg[0][113] = recv_msg[284];
            assign real_msg[0][369] = recv_msg[285];
            assign real_msg[0][241] = recv_msg[286];
            assign real_msg[0][497] = recv_msg[287];
            assign real_msg[0][9] = recv_msg[288];
            assign real_msg[0][265] = recv_msg[289];
            assign real_msg[0][137] = recv_msg[290];
            assign real_msg[0][393] = recv_msg[291];
            assign real_msg[0][73] = recv_msg[292];
            assign real_msg[0][329] = recv_msg[293];
            assign real_msg[0][201] = recv_msg[294];
            assign real_msg[0][457] = recv_msg[295];
            assign real_msg[0][41] = recv_msg[296];
            assign real_msg[0][297] = recv_msg[297];
            assign real_msg[0][169] = recv_msg[298];
            assign real_msg[0][425] = recv_msg[299];
            assign real_msg[0][105] = recv_msg[300];
            assign real_msg[0][361] = recv_msg[301];
            assign real_msg[0][233] = recv_msg[302];
            assign real_msg[0][489] = recv_msg[303];
            assign real_msg[0][25] = recv_msg[304];
            assign real_msg[0][281] = recv_msg[305];
            assign real_msg[0][153] = recv_msg[306];
            assign real_msg[0][409] = recv_msg[307];
            assign real_msg[0][89] = recv_msg[308];
            assign real_msg[0][345] = recv_msg[309];
            assign real_msg[0][217] = recv_msg[310];
            assign real_msg[0][473] = recv_msg[311];
            assign real_msg[0][57] = recv_msg[312];
            assign real_msg[0][313] = recv_msg[313];
            assign real_msg[0][185] = recv_msg[314];
            assign real_msg[0][441] = recv_msg[315];
            assign real_msg[0][121] = recv_msg[316];
            assign real_msg[0][377] = recv_msg[317];
            assign real_msg[0][249] = recv_msg[318];
            assign real_msg[0][505] = recv_msg[319];
            assign real_msg[0][5] = recv_msg[320];
            assign real_msg[0][261] = recv_msg[321];
            assign real_msg[0][133] = recv_msg[322];
            assign real_msg[0][389] = recv_msg[323];
            assign real_msg[0][69] = recv_msg[324];
            assign real_msg[0][325] = recv_msg[325];
            assign real_msg[0][197] = recv_msg[326];
            assign real_msg[0][453] = recv_msg[327];
            assign real_msg[0][37] = recv_msg[328];
            assign real_msg[0][293] = recv_msg[329];
            assign real_msg[0][165] = recv_msg[330];
            assign real_msg[0][421] = recv_msg[331];
            assign real_msg[0][101] = recv_msg[332];
            assign real_msg[0][357] = recv_msg[333];
            assign real_msg[0][229] = recv_msg[334];
            assign real_msg[0][485] = recv_msg[335];
            assign real_msg[0][21] = recv_msg[336];
            assign real_msg[0][277] = recv_msg[337];
            assign real_msg[0][149] = recv_msg[338];
            assign real_msg[0][405] = recv_msg[339];
            assign real_msg[0][85] = recv_msg[340];
            assign real_msg[0][341] = recv_msg[341];
            assign real_msg[0][213] = recv_msg[342];
            assign real_msg[0][469] = recv_msg[343];
            assign real_msg[0][53] = recv_msg[344];
            assign real_msg[0][309] = recv_msg[345];
            assign real_msg[0][181] = recv_msg[346];
            assign real_msg[0][437] = recv_msg[347];
            assign real_msg[0][117] = recv_msg[348];
            assign real_msg[0][373] = recv_msg[349];
            assign real_msg[0][245] = recv_msg[350];
            assign real_msg[0][501] = recv_msg[351];
            assign real_msg[0][13] = recv_msg[352];
            assign real_msg[0][269] = recv_msg[353];
            assign real_msg[0][141] = recv_msg[354];
            assign real_msg[0][397] = recv_msg[355];
            assign real_msg[0][77] = recv_msg[356];
            assign real_msg[0][333] = recv_msg[357];
            assign real_msg[0][205] = recv_msg[358];
            assign real_msg[0][461] = recv_msg[359];
            assign real_msg[0][45] = recv_msg[360];
            assign real_msg[0][301] = recv_msg[361];
            assign real_msg[0][173] = recv_msg[362];
            assign real_msg[0][429] = recv_msg[363];
            assign real_msg[0][109] = recv_msg[364];
            assign real_msg[0][365] = recv_msg[365];
            assign real_msg[0][237] = recv_msg[366];
            assign real_msg[0][493] = recv_msg[367];
            assign real_msg[0][29] = recv_msg[368];
            assign real_msg[0][285] = recv_msg[369];
            assign real_msg[0][157] = recv_msg[370];
            assign real_msg[0][413] = recv_msg[371];
            assign real_msg[0][93] = recv_msg[372];
            assign real_msg[0][349] = recv_msg[373];
            assign real_msg[0][221] = recv_msg[374];
            assign real_msg[0][477] = recv_msg[375];
            assign real_msg[0][61] = recv_msg[376];
            assign real_msg[0][317] = recv_msg[377];
            assign real_msg[0][189] = recv_msg[378];
            assign real_msg[0][445] = recv_msg[379];
            assign real_msg[0][125] = recv_msg[380];
            assign real_msg[0][381] = recv_msg[381];
            assign real_msg[0][253] = recv_msg[382];
            assign real_msg[0][509] = recv_msg[383];
            assign real_msg[0][3] = recv_msg[384];
            assign real_msg[0][259] = recv_msg[385];
            assign real_msg[0][131] = recv_msg[386];
            assign real_msg[0][387] = recv_msg[387];
            assign real_msg[0][67] = recv_msg[388];
            assign real_msg[0][323] = recv_msg[389];
            assign real_msg[0][195] = recv_msg[390];
            assign real_msg[0][451] = recv_msg[391];
            assign real_msg[0][35] = recv_msg[392];
            assign real_msg[0][291] = recv_msg[393];
            assign real_msg[0][163] = recv_msg[394];
            assign real_msg[0][419] = recv_msg[395];
            assign real_msg[0][99] = recv_msg[396];
            assign real_msg[0][355] = recv_msg[397];
            assign real_msg[0][227] = recv_msg[398];
            assign real_msg[0][483] = recv_msg[399];
            assign real_msg[0][19] = recv_msg[400];
            assign real_msg[0][275] = recv_msg[401];
            assign real_msg[0][147] = recv_msg[402];
            assign real_msg[0][403] = recv_msg[403];
            assign real_msg[0][83] = recv_msg[404];
            assign real_msg[0][339] = recv_msg[405];
            assign real_msg[0][211] = recv_msg[406];
            assign real_msg[0][467] = recv_msg[407];
            assign real_msg[0][51] = recv_msg[408];
            assign real_msg[0][307] = recv_msg[409];
            assign real_msg[0][179] = recv_msg[410];
            assign real_msg[0][435] = recv_msg[411];
            assign real_msg[0][115] = recv_msg[412];
            assign real_msg[0][371] = recv_msg[413];
            assign real_msg[0][243] = recv_msg[414];
            assign real_msg[0][499] = recv_msg[415];
            assign real_msg[0][11] = recv_msg[416];
            assign real_msg[0][267] = recv_msg[417];
            assign real_msg[0][139] = recv_msg[418];
            assign real_msg[0][395] = recv_msg[419];
            assign real_msg[0][75] = recv_msg[420];
            assign real_msg[0][331] = recv_msg[421];
            assign real_msg[0][203] = recv_msg[422];
            assign real_msg[0][459] = recv_msg[423];
            assign real_msg[0][43] = recv_msg[424];
            assign real_msg[0][299] = recv_msg[425];
            assign real_msg[0][171] = recv_msg[426];
            assign real_msg[0][427] = recv_msg[427];
            assign real_msg[0][107] = recv_msg[428];
            assign real_msg[0][363] = recv_msg[429];
            assign real_msg[0][235] = recv_msg[430];
            assign real_msg[0][491] = recv_msg[431];
            assign real_msg[0][27] = recv_msg[432];
            assign real_msg[0][283] = recv_msg[433];
            assign real_msg[0][155] = recv_msg[434];
            assign real_msg[0][411] = recv_msg[435];
            assign real_msg[0][91] = recv_msg[436];
            assign real_msg[0][347] = recv_msg[437];
            assign real_msg[0][219] = recv_msg[438];
            assign real_msg[0][475] = recv_msg[439];
            assign real_msg[0][59] = recv_msg[440];
            assign real_msg[0][315] = recv_msg[441];
            assign real_msg[0][187] = recv_msg[442];
            assign real_msg[0][443] = recv_msg[443];
            assign real_msg[0][123] = recv_msg[444];
            assign real_msg[0][379] = recv_msg[445];
            assign real_msg[0][251] = recv_msg[446];
            assign real_msg[0][507] = recv_msg[447];
            assign real_msg[0][7] = recv_msg[448];
            assign real_msg[0][263] = recv_msg[449];
            assign real_msg[0][135] = recv_msg[450];
            assign real_msg[0][391] = recv_msg[451];
            assign real_msg[0][71] = recv_msg[452];
            assign real_msg[0][327] = recv_msg[453];
            assign real_msg[0][199] = recv_msg[454];
            assign real_msg[0][455] = recv_msg[455];
            assign real_msg[0][39] = recv_msg[456];
            assign real_msg[0][295] = recv_msg[457];
            assign real_msg[0][167] = recv_msg[458];
            assign real_msg[0][423] = recv_msg[459];
            assign real_msg[0][103] = recv_msg[460];
            assign real_msg[0][359] = recv_msg[461];
            assign real_msg[0][231] = recv_msg[462];
            assign real_msg[0][487] = recv_msg[463];
            assign real_msg[0][23] = recv_msg[464];
            assign real_msg[0][279] = recv_msg[465];
            assign real_msg[0][151] = recv_msg[466];
            assign real_msg[0][407] = recv_msg[467];
            assign real_msg[0][87] = recv_msg[468];
            assign real_msg[0][343] = recv_msg[469];
            assign real_msg[0][215] = recv_msg[470];
            assign real_msg[0][471] = recv_msg[471];
            assign real_msg[0][55] = recv_msg[472];
            assign real_msg[0][311] = recv_msg[473];
            assign real_msg[0][183] = recv_msg[474];
            assign real_msg[0][439] = recv_msg[475];
            assign real_msg[0][119] = recv_msg[476];
            assign real_msg[0][375] = recv_msg[477];
            assign real_msg[0][247] = recv_msg[478];
            assign real_msg[0][503] = recv_msg[479];
            assign real_msg[0][15] = recv_msg[480];
            assign real_msg[0][271] = recv_msg[481];
            assign real_msg[0][143] = recv_msg[482];
            assign real_msg[0][399] = recv_msg[483];
            assign real_msg[0][79] = recv_msg[484];
            assign real_msg[0][335] = recv_msg[485];
            assign real_msg[0][207] = recv_msg[486];
            assign real_msg[0][463] = recv_msg[487];
            assign real_msg[0][47] = recv_msg[488];
            assign real_msg[0][303] = recv_msg[489];
            assign real_msg[0][175] = recv_msg[490];
            assign real_msg[0][431] = recv_msg[491];
            assign real_msg[0][111] = recv_msg[492];
            assign real_msg[0][367] = recv_msg[493];
            assign real_msg[0][239] = recv_msg[494];
            assign real_msg[0][495] = recv_msg[495];
            assign real_msg[0][31] = recv_msg[496];
            assign real_msg[0][287] = recv_msg[497];
            assign real_msg[0][159] = recv_msg[498];
            assign real_msg[0][415] = recv_msg[499];
            assign real_msg[0][95] = recv_msg[500];
            assign real_msg[0][351] = recv_msg[501];
            assign real_msg[0][223] = recv_msg[502];
            assign real_msg[0][479] = recv_msg[503];
            assign real_msg[0][63] = recv_msg[504];
            assign real_msg[0][319] = recv_msg[505];
            assign real_msg[0][191] = recv_msg[506];
            assign real_msg[0][447] = recv_msg[507];
            assign real_msg[0][127] = recv_msg[508];
            assign real_msg[0][383] = recv_msg[509];
            assign real_msg[0][255] = recv_msg[510];
            assign real_msg[0][511] = recv_msg[511];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_512VRTL SineWave (.sine_wave_out(sine_wave_out));
        end else if(N_SAMPLES == 256) begin
           assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][128] = recv_msg[1];
            assign real_msg[0][64] = recv_msg[2];
            assign real_msg[0][192] = recv_msg[3];
            assign real_msg[0][32] = recv_msg[4];
            assign real_msg[0][160] = recv_msg[5];
            assign real_msg[0][96] = recv_msg[6];
            assign real_msg[0][224] = recv_msg[7];
            assign real_msg[0][16] = recv_msg[8];
            assign real_msg[0][144] = recv_msg[9];
            assign real_msg[0][80] = recv_msg[10];
            assign real_msg[0][208] = recv_msg[11];
            assign real_msg[0][48] = recv_msg[12];
            assign real_msg[0][176] = recv_msg[13];
            assign real_msg[0][112] = recv_msg[14];
            assign real_msg[0][240] = recv_msg[15];
            assign real_msg[0][8] = recv_msg[16];
            assign real_msg[0][136] = recv_msg[17];
            assign real_msg[0][72] = recv_msg[18];
            assign real_msg[0][200] = recv_msg[19];
            assign real_msg[0][40] = recv_msg[20];
            assign real_msg[0][168] = recv_msg[21];
            assign real_msg[0][104] = recv_msg[22];
            assign real_msg[0][232] = recv_msg[23];
            assign real_msg[0][24] = recv_msg[24];
            assign real_msg[0][152] = recv_msg[25];
            assign real_msg[0][88] = recv_msg[26];
            assign real_msg[0][216] = recv_msg[27];
            assign real_msg[0][56] = recv_msg[28];
            assign real_msg[0][184] = recv_msg[29];
            assign real_msg[0][120] = recv_msg[30];
            assign real_msg[0][248] = recv_msg[31];
            assign real_msg[0][4] = recv_msg[32];
            assign real_msg[0][132] = recv_msg[33];
            assign real_msg[0][68] = recv_msg[34];
            assign real_msg[0][196] = recv_msg[35];
            assign real_msg[0][36] = recv_msg[36];
            assign real_msg[0][164] = recv_msg[37];
            assign real_msg[0][100] = recv_msg[38];
            assign real_msg[0][228] = recv_msg[39];
            assign real_msg[0][20] = recv_msg[40];
            assign real_msg[0][148] = recv_msg[41];
            assign real_msg[0][84] = recv_msg[42];
            assign real_msg[0][212] = recv_msg[43];
            assign real_msg[0][52] = recv_msg[44];
            assign real_msg[0][180] = recv_msg[45];
            assign real_msg[0][116] = recv_msg[46];
            assign real_msg[0][244] = recv_msg[47];
            assign real_msg[0][12] = recv_msg[48];
            assign real_msg[0][140] = recv_msg[49];
            assign real_msg[0][76] = recv_msg[50];
            assign real_msg[0][204] = recv_msg[51];
            assign real_msg[0][44] = recv_msg[52];
            assign real_msg[0][172] = recv_msg[53];
            assign real_msg[0][108] = recv_msg[54];
            assign real_msg[0][236] = recv_msg[55];
            assign real_msg[0][28] = recv_msg[56];
            assign real_msg[0][156] = recv_msg[57];
            assign real_msg[0][92] = recv_msg[58];
            assign real_msg[0][220] = recv_msg[59];
            assign real_msg[0][60] = recv_msg[60];
            assign real_msg[0][188] = recv_msg[61];
            assign real_msg[0][124] = recv_msg[62];
            assign real_msg[0][252] = recv_msg[63];
            assign real_msg[0][2] = recv_msg[64];
            assign real_msg[0][130] = recv_msg[65];
            assign real_msg[0][66] = recv_msg[66];
            assign real_msg[0][194] = recv_msg[67];
            assign real_msg[0][34] = recv_msg[68];
            assign real_msg[0][162] = recv_msg[69];
            assign real_msg[0][98] = recv_msg[70];
            assign real_msg[0][226] = recv_msg[71];
            assign real_msg[0][18] = recv_msg[72];
            assign real_msg[0][146] = recv_msg[73];
            assign real_msg[0][82] = recv_msg[74];
            assign real_msg[0][210] = recv_msg[75];
            assign real_msg[0][50] = recv_msg[76];
            assign real_msg[0][178] = recv_msg[77];
            assign real_msg[0][114] = recv_msg[78];
            assign real_msg[0][242] = recv_msg[79];
            assign real_msg[0][10] = recv_msg[80];
            assign real_msg[0][138] = recv_msg[81];
            assign real_msg[0][74] = recv_msg[82];
            assign real_msg[0][202] = recv_msg[83];
            assign real_msg[0][42] = recv_msg[84];
            assign real_msg[0][170] = recv_msg[85];
            assign real_msg[0][106] = recv_msg[86];
            assign real_msg[0][234] = recv_msg[87];
            assign real_msg[0][26] = recv_msg[88];
            assign real_msg[0][154] = recv_msg[89];
            assign real_msg[0][90] = recv_msg[90];
            assign real_msg[0][218] = recv_msg[91];
            assign real_msg[0][58] = recv_msg[92];
            assign real_msg[0][186] = recv_msg[93];
            assign real_msg[0][122] = recv_msg[94];
            assign real_msg[0][250] = recv_msg[95];
            assign real_msg[0][6] = recv_msg[96];
            assign real_msg[0][134] = recv_msg[97];
            assign real_msg[0][70] = recv_msg[98];
            assign real_msg[0][198] = recv_msg[99];
            assign real_msg[0][38] = recv_msg[100];
            assign real_msg[0][166] = recv_msg[101];
            assign real_msg[0][102] = recv_msg[102];
            assign real_msg[0][230] = recv_msg[103];
            assign real_msg[0][22] = recv_msg[104];
            assign real_msg[0][150] = recv_msg[105];
            assign real_msg[0][86] = recv_msg[106];
            assign real_msg[0][214] = recv_msg[107];
            assign real_msg[0][54] = recv_msg[108];
            assign real_msg[0][182] = recv_msg[109];
            assign real_msg[0][118] = recv_msg[110];
            assign real_msg[0][246] = recv_msg[111];
            assign real_msg[0][14] = recv_msg[112];
            assign real_msg[0][142] = recv_msg[113];
            assign real_msg[0][78] = recv_msg[114];
            assign real_msg[0][206] = recv_msg[115];
            assign real_msg[0][46] = recv_msg[116];
            assign real_msg[0][174] = recv_msg[117];
            assign real_msg[0][110] = recv_msg[118];
            assign real_msg[0][238] = recv_msg[119];
            assign real_msg[0][30] = recv_msg[120];
            assign real_msg[0][158] = recv_msg[121];
            assign real_msg[0][94] = recv_msg[122];
            assign real_msg[0][222] = recv_msg[123];
            assign real_msg[0][62] = recv_msg[124];
            assign real_msg[0][190] = recv_msg[125];
            assign real_msg[0][126] = recv_msg[126];
            assign real_msg[0][254] = recv_msg[127];
            assign real_msg[0][1] = recv_msg[128];
            assign real_msg[0][129] = recv_msg[129];
            assign real_msg[0][65] = recv_msg[130];
            assign real_msg[0][193] = recv_msg[131];
            assign real_msg[0][33] = recv_msg[132];
            assign real_msg[0][161] = recv_msg[133];
            assign real_msg[0][97] = recv_msg[134];
            assign real_msg[0][225] = recv_msg[135];
            assign real_msg[0][17] = recv_msg[136];
            assign real_msg[0][145] = recv_msg[137];
            assign real_msg[0][81] = recv_msg[138];
            assign real_msg[0][209] = recv_msg[139];
            assign real_msg[0][49] = recv_msg[140];
            assign real_msg[0][177] = recv_msg[141];
            assign real_msg[0][113] = recv_msg[142];
            assign real_msg[0][241] = recv_msg[143];
            assign real_msg[0][9] = recv_msg[144];
            assign real_msg[0][137] = recv_msg[145];
            assign real_msg[0][73] = recv_msg[146];
            assign real_msg[0][201] = recv_msg[147];
            assign real_msg[0][41] = recv_msg[148];
            assign real_msg[0][169] = recv_msg[149];
            assign real_msg[0][105] = recv_msg[150];
            assign real_msg[0][233] = recv_msg[151];
            assign real_msg[0][25] = recv_msg[152];
            assign real_msg[0][153] = recv_msg[153];
            assign real_msg[0][89] = recv_msg[154];
            assign real_msg[0][217] = recv_msg[155];
            assign real_msg[0][57] = recv_msg[156];
            assign real_msg[0][185] = recv_msg[157];
            assign real_msg[0][121] = recv_msg[158];
            assign real_msg[0][249] = recv_msg[159];
            assign real_msg[0][5] = recv_msg[160];
            assign real_msg[0][133] = recv_msg[161];
            assign real_msg[0][69] = recv_msg[162];
            assign real_msg[0][197] = recv_msg[163];
            assign real_msg[0][37] = recv_msg[164];
            assign real_msg[0][165] = recv_msg[165];
            assign real_msg[0][101] = recv_msg[166];
            assign real_msg[0][229] = recv_msg[167];
            assign real_msg[0][21] = recv_msg[168];
            assign real_msg[0][149] = recv_msg[169];
            assign real_msg[0][85] = recv_msg[170];
            assign real_msg[0][213] = recv_msg[171];
            assign real_msg[0][53] = recv_msg[172];
            assign real_msg[0][181] = recv_msg[173];
            assign real_msg[0][117] = recv_msg[174];
            assign real_msg[0][245] = recv_msg[175];
            assign real_msg[0][13] = recv_msg[176];
            assign real_msg[0][141] = recv_msg[177];
            assign real_msg[0][77] = recv_msg[178];
            assign real_msg[0][205] = recv_msg[179];
            assign real_msg[0][45] = recv_msg[180];
            assign real_msg[0][173] = recv_msg[181];
            assign real_msg[0][109] = recv_msg[182];
            assign real_msg[0][237] = recv_msg[183];
            assign real_msg[0][29] = recv_msg[184];
            assign real_msg[0][157] = recv_msg[185];
            assign real_msg[0][93] = recv_msg[186];
            assign real_msg[0][221] = recv_msg[187];
            assign real_msg[0][61] = recv_msg[188];
            assign real_msg[0][189] = recv_msg[189];
            assign real_msg[0][125] = recv_msg[190];
            assign real_msg[0][253] = recv_msg[191];
            assign real_msg[0][3] = recv_msg[192];
            assign real_msg[0][131] = recv_msg[193];
            assign real_msg[0][67] = recv_msg[194];
            assign real_msg[0][195] = recv_msg[195];
            assign real_msg[0][35] = recv_msg[196];
            assign real_msg[0][163] = recv_msg[197];
            assign real_msg[0][99] = recv_msg[198];
            assign real_msg[0][227] = recv_msg[199];
            assign real_msg[0][19] = recv_msg[200];
            assign real_msg[0][147] = recv_msg[201];
            assign real_msg[0][83] = recv_msg[202];
            assign real_msg[0][211] = recv_msg[203];
            assign real_msg[0][51] = recv_msg[204];
            assign real_msg[0][179] = recv_msg[205];
            assign real_msg[0][115] = recv_msg[206];
            assign real_msg[0][243] = recv_msg[207];
            assign real_msg[0][11] = recv_msg[208];
            assign real_msg[0][139] = recv_msg[209];
            assign real_msg[0][75] = recv_msg[210];
            assign real_msg[0][203] = recv_msg[211];
            assign real_msg[0][43] = recv_msg[212];
            assign real_msg[0][171] = recv_msg[213];
            assign real_msg[0][107] = recv_msg[214];
            assign real_msg[0][235] = recv_msg[215];
            assign real_msg[0][27] = recv_msg[216];
            assign real_msg[0][155] = recv_msg[217];
            assign real_msg[0][91] = recv_msg[218];
            assign real_msg[0][219] = recv_msg[219];
            assign real_msg[0][59] = recv_msg[220];
            assign real_msg[0][187] = recv_msg[221];
            assign real_msg[0][123] = recv_msg[222];
            assign real_msg[0][251] = recv_msg[223];
            assign real_msg[0][7] = recv_msg[224];
            assign real_msg[0][135] = recv_msg[225];
            assign real_msg[0][71] = recv_msg[226];
            assign real_msg[0][199] = recv_msg[227];
            assign real_msg[0][39] = recv_msg[228];
            assign real_msg[0][167] = recv_msg[229];
            assign real_msg[0][103] = recv_msg[230];
            assign real_msg[0][231] = recv_msg[231];
            assign real_msg[0][23] = recv_msg[232];
            assign real_msg[0][151] = recv_msg[233];
            assign real_msg[0][87] = recv_msg[234];
            assign real_msg[0][215] = recv_msg[235];
            assign real_msg[0][55] = recv_msg[236];
            assign real_msg[0][183] = recv_msg[237];
            assign real_msg[0][119] = recv_msg[238];
            assign real_msg[0][247] = recv_msg[239];
            assign real_msg[0][15] = recv_msg[240];
            assign real_msg[0][143] = recv_msg[241];
            assign real_msg[0][79] = recv_msg[242];
            assign real_msg[0][207] = recv_msg[243];
            assign real_msg[0][47] = recv_msg[244];
            assign real_msg[0][175] = recv_msg[245];
            assign real_msg[0][111] = recv_msg[246];
            assign real_msg[0][239] = recv_msg[247];
            assign real_msg[0][31] = recv_msg[248];
            assign real_msg[0][159] = recv_msg[249];
            assign real_msg[0][95] = recv_msg[250];
            assign real_msg[0][223] = recv_msg[251];
            assign real_msg[0][63] = recv_msg[252];
            assign real_msg[0][191] = recv_msg[253];
            assign real_msg[0][127] = recv_msg[254];
            assign real_msg[0][255] = recv_msg[255];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_256VRTL SineWave (.sine_wave_out(sine_wave_out));
        
        end else if(N_SAMPLES == 128) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][64] = recv_msg[1];
            assign real_msg[0][32] = recv_msg[2];
            assign real_msg[0][96] = recv_msg[3];
            assign real_msg[0][16] = recv_msg[4];
            assign real_msg[0][80] = recv_msg[5];
            assign real_msg[0][48] = recv_msg[6];
            assign real_msg[0][112] = recv_msg[7];
            assign real_msg[0][8] = recv_msg[8];
            assign real_msg[0][72] = recv_msg[9];
            assign real_msg[0][40] = recv_msg[10];
            assign real_msg[0][104] = recv_msg[11];
            assign real_msg[0][24] = recv_msg[12];
            assign real_msg[0][88] = recv_msg[13];
            assign real_msg[0][56] = recv_msg[14];
            assign real_msg[0][120] = recv_msg[15];
            assign real_msg[0][4] = recv_msg[16];
            assign real_msg[0][68] = recv_msg[17];
            assign real_msg[0][36] = recv_msg[18];
            assign real_msg[0][100] = recv_msg[19];
            assign real_msg[0][20] = recv_msg[20];
            assign real_msg[0][84] = recv_msg[21];
            assign real_msg[0][52] = recv_msg[22];
            assign real_msg[0][116] = recv_msg[23];
            assign real_msg[0][12] = recv_msg[24];
            assign real_msg[0][76] = recv_msg[25];
            assign real_msg[0][44] = recv_msg[26];
            assign real_msg[0][108] = recv_msg[27];
            assign real_msg[0][28] = recv_msg[28];
            assign real_msg[0][92] = recv_msg[29];
            assign real_msg[0][60] = recv_msg[30];
            assign real_msg[0][124] = recv_msg[31];
            assign real_msg[0][2] = recv_msg[32];
            assign real_msg[0][66] = recv_msg[33];
            assign real_msg[0][34] = recv_msg[34];
            assign real_msg[0][98] = recv_msg[35];
            assign real_msg[0][18] = recv_msg[36];
            assign real_msg[0][82] = recv_msg[37];
            assign real_msg[0][50] = recv_msg[38];
            assign real_msg[0][114] = recv_msg[39];
            assign real_msg[0][10] = recv_msg[40];
            assign real_msg[0][74] = recv_msg[41];
            assign real_msg[0][42] = recv_msg[42];
            assign real_msg[0][106] = recv_msg[43];
            assign real_msg[0][26] = recv_msg[44];
            assign real_msg[0][90] = recv_msg[45];
            assign real_msg[0][58] = recv_msg[46];
            assign real_msg[0][122] = recv_msg[47];
            assign real_msg[0][6] = recv_msg[48];
            assign real_msg[0][70] = recv_msg[49];
            assign real_msg[0][38] = recv_msg[50];
            assign real_msg[0][102] = recv_msg[51];
            assign real_msg[0][22] = recv_msg[52];
            assign real_msg[0][86] = recv_msg[53];
            assign real_msg[0][54] = recv_msg[54];
            assign real_msg[0][118] = recv_msg[55];
            assign real_msg[0][14] = recv_msg[56];
            assign real_msg[0][78] = recv_msg[57];
            assign real_msg[0][46] = recv_msg[58];
            assign real_msg[0][110] = recv_msg[59];
            assign real_msg[0][30] = recv_msg[60];
            assign real_msg[0][94] = recv_msg[61];
            assign real_msg[0][62] = recv_msg[62];
            assign real_msg[0][126] = recv_msg[63];
            assign real_msg[0][1] = recv_msg[64];
            assign real_msg[0][65] = recv_msg[65];
            assign real_msg[0][33] = recv_msg[66];
            assign real_msg[0][97] = recv_msg[67];
            assign real_msg[0][17] = recv_msg[68];
            assign real_msg[0][81] = recv_msg[69];
            assign real_msg[0][49] = recv_msg[70];
            assign real_msg[0][113] = recv_msg[71];
            assign real_msg[0][9] = recv_msg[72];
            assign real_msg[0][73] = recv_msg[73];
            assign real_msg[0][41] = recv_msg[74];
            assign real_msg[0][105] = recv_msg[75];
            assign real_msg[0][25] = recv_msg[76];
            assign real_msg[0][89] = recv_msg[77];
            assign real_msg[0][57] = recv_msg[78];
            assign real_msg[0][121] = recv_msg[79];
            assign real_msg[0][5] = recv_msg[80];
            assign real_msg[0][69] = recv_msg[81];
            assign real_msg[0][37] = recv_msg[82];
            assign real_msg[0][101] = recv_msg[83];
            assign real_msg[0][21] = recv_msg[84];
            assign real_msg[0][85] = recv_msg[85];
            assign real_msg[0][53] = recv_msg[86];
            assign real_msg[0][117] = recv_msg[87];
            assign real_msg[0][13] = recv_msg[88];
            assign real_msg[0][77] = recv_msg[89];
            assign real_msg[0][45] = recv_msg[90];
            assign real_msg[0][109] = recv_msg[91];
            assign real_msg[0][29] = recv_msg[92];
            assign real_msg[0][93] = recv_msg[93];
            assign real_msg[0][61] = recv_msg[94];
            assign real_msg[0][125] = recv_msg[95];
            assign real_msg[0][3] = recv_msg[96];
            assign real_msg[0][67] = recv_msg[97];
            assign real_msg[0][35] = recv_msg[98];
            assign real_msg[0][99] = recv_msg[99];
            assign real_msg[0][19] = recv_msg[100];
            assign real_msg[0][83] = recv_msg[101];
            assign real_msg[0][51] = recv_msg[102];
            assign real_msg[0][115] = recv_msg[103];
            assign real_msg[0][11] = recv_msg[104];
            assign real_msg[0][75] = recv_msg[105];
            assign real_msg[0][43] = recv_msg[106];
            assign real_msg[0][107] = recv_msg[107];
            assign real_msg[0][27] = recv_msg[108];
            assign real_msg[0][91] = recv_msg[109];
            assign real_msg[0][59] = recv_msg[110];
            assign real_msg[0][123] = recv_msg[111];
            assign real_msg[0][7] = recv_msg[112];
            assign real_msg[0][71] = recv_msg[113];
            assign real_msg[0][39] = recv_msg[114];
            assign real_msg[0][103] = recv_msg[115];
            assign real_msg[0][23] = recv_msg[116];
            assign real_msg[0][87] = recv_msg[117];
            assign real_msg[0][55] = recv_msg[118];
            assign real_msg[0][119] = recv_msg[119];
            assign real_msg[0][15] = recv_msg[120];
            assign real_msg[0][79] = recv_msg[121];
            assign real_msg[0][47] = recv_msg[122];
            assign real_msg[0][111] = recv_msg[123];
            assign real_msg[0][31] = recv_msg[124];
            assign real_msg[0][95] = recv_msg[125];
            assign real_msg[0][63] = recv_msg[126];
            assign real_msg[0][127] = recv_msg[127];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_128VRTL SineWave (.sine_wave_out(sine_wave_out));
        end else if(N_SAMPLES == 64) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][32] = recv_msg[1];
            assign real_msg[0][16] = recv_msg[2];
            assign real_msg[0][48] = recv_msg[3];
            assign real_msg[0][8] = recv_msg[4];
            assign real_msg[0][40] = recv_msg[5];
            assign real_msg[0][24] = recv_msg[6];
            assign real_msg[0][56] = recv_msg[7];
            assign real_msg[0][4] = recv_msg[8];
            assign real_msg[0][36] = recv_msg[9];
            assign real_msg[0][20] = recv_msg[10];
            assign real_msg[0][52] = recv_msg[11];
            assign real_msg[0][12] = recv_msg[12];
            assign real_msg[0][44] = recv_msg[13];
            assign real_msg[0][28] = recv_msg[14];
            assign real_msg[0][60] = recv_msg[15];
            assign real_msg[0][2] = recv_msg[16];
            assign real_msg[0][34] = recv_msg[17];
            assign real_msg[0][18] = recv_msg[18];
            assign real_msg[0][50] = recv_msg[19];
            assign real_msg[0][10] = recv_msg[20];
            assign real_msg[0][42] = recv_msg[21];
            assign real_msg[0][26] = recv_msg[22];
            assign real_msg[0][58] = recv_msg[23];
            assign real_msg[0][6] = recv_msg[24];
            assign real_msg[0][38] = recv_msg[25];
            assign real_msg[0][22] = recv_msg[26];
            assign real_msg[0][54] = recv_msg[27];
            assign real_msg[0][14] = recv_msg[28];
            assign real_msg[0][46] = recv_msg[29];
            assign real_msg[0][30] = recv_msg[30];
            assign real_msg[0][62] = recv_msg[31];
            assign real_msg[0][1] = recv_msg[32];
            assign real_msg[0][33] = recv_msg[33];
            assign real_msg[0][17] = recv_msg[34];
            assign real_msg[0][49] = recv_msg[35];
            assign real_msg[0][9] = recv_msg[36];
            assign real_msg[0][41] = recv_msg[37];
            assign real_msg[0][25] = recv_msg[38];
            assign real_msg[0][57] = recv_msg[39];
            assign real_msg[0][5] = recv_msg[40];
            assign real_msg[0][37] = recv_msg[41];
            assign real_msg[0][21] = recv_msg[42];
            assign real_msg[0][53] = recv_msg[43];
            assign real_msg[0][13] = recv_msg[44];
            assign real_msg[0][45] = recv_msg[45];
            assign real_msg[0][29] = recv_msg[46];
            assign real_msg[0][61] = recv_msg[47];
            assign real_msg[0][3] = recv_msg[48];
            assign real_msg[0][35] = recv_msg[49];
            assign real_msg[0][19] = recv_msg[50];
            assign real_msg[0][51] = recv_msg[51];
            assign real_msg[0][11] = recv_msg[52];
            assign real_msg[0][43] = recv_msg[53];
            assign real_msg[0][27] = recv_msg[54];
            assign real_msg[0][59] = recv_msg[55];
            assign real_msg[0][7] = recv_msg[56];
            assign real_msg[0][39] = recv_msg[57];
            assign real_msg[0][23] = recv_msg[58];
            assign real_msg[0][55] = recv_msg[59];
            assign real_msg[0][15] = recv_msg[60];
            assign real_msg[0][47] = recv_msg[61];
            assign real_msg[0][31] = recv_msg[62];
            assign real_msg[0][63] = recv_msg[63];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_64VRTL SineWave (.sine_wave_out(sine_wave_out));

        end else if(N_SAMPLES == 32) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][16] = recv_msg[1];
            assign real_msg[0][8] = recv_msg[2];
            assign real_msg[0][24] = recv_msg[3];
            assign real_msg[0][4] = recv_msg[4];
            assign real_msg[0][20] = recv_msg[5];
            assign real_msg[0][12] = recv_msg[6];
            assign real_msg[0][28] = recv_msg[7];
            assign real_msg[0][2] = recv_msg[8];
            assign real_msg[0][18] = recv_msg[9];
            assign real_msg[0][10] = recv_msg[10];
            assign real_msg[0][26] = recv_msg[11];
            assign real_msg[0][6] = recv_msg[12];
            assign real_msg[0][22] = recv_msg[13];
            assign real_msg[0][14] = recv_msg[14];
            assign real_msg[0][30] = recv_msg[15];
            assign real_msg[0][1] = recv_msg[16];
            assign real_msg[0][17] = recv_msg[17];
            assign real_msg[0][9] = recv_msg[18];
            assign real_msg[0][25] = recv_msg[19];
            assign real_msg[0][5] = recv_msg[20];
            assign real_msg[0][21] = recv_msg[21];
            assign real_msg[0][13] = recv_msg[22];
            assign real_msg[0][29] = recv_msg[23];
            assign real_msg[0][3] = recv_msg[24];
            assign real_msg[0][19] = recv_msg[25];
            assign real_msg[0][11] = recv_msg[26];
            assign real_msg[0][27] = recv_msg[27];
            assign real_msg[0][7] = recv_msg[28];
            assign real_msg[0][23] = recv_msg[29];
            assign real_msg[0][15] = recv_msg[30];
            assign real_msg[0][31] = recv_msg[31];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_32VRTL SineWave (.sine_wave_out(sine_wave_out));

        end else if(N_SAMPLES == 16) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][8] = recv_msg[1];
            assign real_msg[0][4] = recv_msg[2];
            assign real_msg[0][12] = recv_msg[3];
            assign real_msg[0][2] = recv_msg[4];
            assign real_msg[0][10] = recv_msg[5];
            assign real_msg[0][6] = recv_msg[6];
            assign real_msg[0][14] = recv_msg[7];
            assign real_msg[0][1] = recv_msg[8];
            assign real_msg[0][9] = recv_msg[9];
            assign real_msg[0][5] = recv_msg[10];
            assign real_msg[0][13] = recv_msg[11];
            assign real_msg[0][3] = recv_msg[12];
            assign real_msg[0][11] = recv_msg[13];
            assign real_msg[0][7] = recv_msg[14];
            assign real_msg[0][15] = recv_msg[15];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_16VRTL SineWave (.sine_wave_out(sine_wave_out));

        end else if(N_SAMPLES == 8) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][4] = recv_msg[1];
            assign real_msg[0][2] = recv_msg[2];
            assign real_msg[0][6] = recv_msg[3];
            assign real_msg[0][1] = recv_msg[4];
            assign real_msg[0][5] = recv_msg[5];
            assign real_msg[0][3] = recv_msg[6];
            assign real_msg[0][7] = recv_msg[7];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_8VRTL SineWave (.sine_wave_out(sine_wave_out));

        end else if(N_SAMPLES == 4) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][2] = recv_msg[1];
            assign real_msg[0][1] = recv_msg[2];
            assign real_msg[0][3] = recv_msg[3];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_4VRTL SineWave (.sine_wave_out(sine_wave_out));
			
        end else if(N_SAMPLES == 2) begin
            assign real_msg[0][0] = recv_msg[0];
            assign real_msg[0][1] = recv_msg[1];
            SineWave__BIT_WIDTH_32__DECIMAL_POINT_16__SIZE_FFT_2VRTL SineWave (.sine_wave_out(sine_wave_out));

        end
    endgenerate

    
    
    generate
        genvar i;
        genvar b;
        for( i = 0; i < $clog2(N_SAMPLES); i++ ) begin
            FFT_StageVRTL #(.BIT_WIDTH(BIT_WIDTH), .DECIMAL_PT(DECIMAL_PT), .N_SAMPLES(N_SAMPLES), .STAGE_FFT(i)) fft_stage ( 
                .recv_msg_real(real_msg   [i]),
                .recv_msg_imag(complex_msg[i]),
                .recv_val     (val_in     [i]),
                .recv_rdy     (rdy_in     [i]),
        
                .send_msg_real(real_msg   [i + 1]),
                .send_msg_imag(complex_msg[i + 1]),
                .send_val     (val_in     [i + 1]),
                .send_rdy     (rdy_in     [i + 1]),

                .sine_wave_out(sine_wave_out),

                .reset        (reset),
                .clk          (clk)
                );
        end
    endgenerate

    always @(*) begin
        int i;
        for(i = 0; i < N_SAMPLES; i++) begin

            send_msg[i] = real_msg[$clog2(N_SAMPLES)][i];

        end
    end
    

endmodule

`endif